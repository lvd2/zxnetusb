// ZXiznet project
// (c) NedoPC 2012
//
// mapping of wiznet address space

module wizmap
(
);



endmodule

