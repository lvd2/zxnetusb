// ZXiznet project
// (c) NedoPC 2012
//
// all zx-bus functions

module zbus
(
);


endmodule

